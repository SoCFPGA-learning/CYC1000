module constant(
    output wire const
);
   
assign const = 1'b1;
    
endmodule
